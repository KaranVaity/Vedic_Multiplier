** Profile: "SCHEMATIC1-test"  [ C:\Users\Karan\Documents\PSpice\VLSI\vlsi-schematic1-test.sim ] 

** Creating circuit file "vlsi-schematic1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad 9.1\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ns 0 1ns 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\vlsi-SCHEMATIC1.net" 


.END
