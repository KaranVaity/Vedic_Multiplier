** Profile: "MAIN-test2"  [ C:\Users\Karan\Documents\PSpice\VLSI\vlsi-main-test2.sim ] 

** Creating circuit file "vlsi-main-test2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.STMLIB ".\VLSI.stl" 
* From [PSPICE NETLIST] section of C:\Program Files\Orcad 9.1\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 40ms 0 0.1ms 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\vlsi-MAIN.net" 


.END
