** Profile: "MAIN-test4"  [ C:\Users\Karan\Documents\PSpice\VLSI\vlsi-MAIN-test4.sim ] 

** Creating circuit file "vlsi-MAIN-test4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.STMLIB ".\VLSI.stl" 
* From [PSPICE NETLIST] section of C:\Program Files\Orcad 9.1\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\vlsi-MAIN.net" 


.END
